module avg (
  input logic rst_ni,
  input logic clk_i,
  input logic data_i,
  output logic data_o
);



endmodule