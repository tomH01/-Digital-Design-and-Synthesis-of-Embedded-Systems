module and_gate (
    input logic a, b,
    output o
);
    assign o = a & b;
endmodule    
